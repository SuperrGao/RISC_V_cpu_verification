`ifndef MY_SCOREBOARD__SV
`define MY_SCOREBOARD__SV
class my_scoreboard extends uvm_scoreboard;
	my_transaction  expect_queue[$];
	uvm_blocking_get_port #(my_transaction)  exp_port;
	uvm_blocking_get_port #(my_transaction)  act_port;
	`uvm_component_utils(my_scoreboard)
	
	extern function new(string name, uvm_component parent = null);
	extern virtual function void build_phase(uvm_phase phase);
	extern virtual task main_phase(uvm_phase phase);
endclass 

function my_scoreboard::new(string name, uvm_component parent = null);
	super.new(name, parent);
endfunction 

function void my_scoreboard::build_phase(uvm_phase phase);
	super.build_phase(phase);
	exp_port = new("exp_port", this);
	act_port = new("act_port", this);
endfunction 

task my_scoreboard::main_phase(uvm_phase phase);
	my_transaction  get_expect,  get_actual, tmp_tran;
	bit result;
	super.main_phase(phase);
	fork 
		while (1) begin
			exp_port.get(get_expect);
			`uvm_info("my_scoreboard", "get one transaction model", UVM_LOW)
			expect_queue.push_back(get_expect);
		end
		while (1) begin
			act_port.get(get_actual);
			#1
			`uvm_info("my_scoreboard", "get one transaction from dut", UVM_LOW)
			if(expect_queue.size() > 0) begin
				tmp_tran = expect_queue.pop_front();
				result =    (get_actual.s0_addr   == tmp_tran.s0_addr)   && (get_actual.s1_addr   == tmp_tran.s1_addr)   &&
							(get_actual.s2_addr   == tmp_tran.s2_addr)   && (get_actual.s3_addr   == tmp_tran.s3_addr)   &&
							(get_actual.s4_addr   == tmp_tran.s4_addr)   && (get_actual.s5_addr   == tmp_tran.s5_addr)   &&
							(get_actual.m0_data_o == tmp_tran.m0_data_o) && (get_actual.m1_data_o == tmp_tran.m1_data_o) &&
							(get_actual.m2_data_o == tmp_tran.m2_data_o) && (get_actual.m3_data_o == tmp_tran.m3_data_o) &&
							(get_actual.s0_data_o == tmp_tran.s0_data_o) && (get_actual.s1_data_o == tmp_tran.s1_data_o) &&
							(get_actual.s2_data_o == tmp_tran.s2_data_o) && (get_actual.s3_data_o == tmp_tran.s3_data_o) &&
							(get_actual.s4_data_o == tmp_tran.s4_data_o) && (get_actual.s5_data_o == tmp_tran.s5_data_o);
							/*get_actual.hold_flag === tmp_tran.hold_flag*/

				if(result) begin 
					`uvm_info("my_scoreboard", "Compare SUCCESSFULLY", UVM_LOW);
					$display("the expect pkt is");
					tmp_tran.print();
					$display("the actual pkt is");
					get_actual.print();
				end
				else begin
					`uvm_error("my_scoreboard", "Compare FAILED");
					$display("the expect pkt is");
					tmp_tran.print();
					$display("the actual pkt is");
					get_actual.print();
				end
			end
			else begin
				`uvm_error("my_scoreboard", "Received from DUT, while Expect Queue is empty");
				$display("the unexpected pkt is");
				get_actual.print();
			end 
		end
	join
endtask
`endif
